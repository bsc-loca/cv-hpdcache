/*
 *  Copyright 2023 CEA*
 *  *Commissariat a l'Energie Atomique et aux Energies Alternatives (CEA)
 *
 *  SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 *
 *  Licensed under the Solderpad Hardware License v 2.1 (the “License”); you
 *  may not use this file except in compliance with the License, or, at your
 *  option, the Apache License version 2.0. You may obtain a copy of the
 *  License at
 *
 *  https://solderpad.org/licenses/SHL-2.1/
 *
 *  Unless required by applicable law or agreed to in writing, any work
 *  distributed under the License is distributed on an “AS IS” BASIS, WITHOUT
 *  WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
 *  License for the specific language governing permissions and limitations
 *  under the License.
 */
/*
 *  Authors       : Cesar Fuguet
 *  Creation Date : March, 2020
 *  Description   : Wrapper for Behavioral SRAM macros
 *  History       :
 */
module hpdcache_sram
#(
    parameter int unsigned ADDR_SIZE = 0,
    parameter int unsigned DATA_SIZE = 0,
    parameter int unsigned DEPTH = 2**ADDR_SIZE
)
(
    `ifdef INTEL_PHYSICAL_MEM_CTRL
    input  logic [27:0]           uhdusplr_mem_ctrl,
    `endif
    input  logic                  clk,
    input  logic                  rst_n,
    input  logic                  cs,
    input  logic                  we,
    input  logic [ADDR_SIZE-1:0]  addr,
    input  logic [DATA_SIZE-1:0]  wdata,
    output logic [DATA_SIZE-1:0]  rdata
);

    sp_ram #(
        .ADDR_WIDTH(ADDR_SIZE),
        .DATA_WIDTH(DATA_SIZE),
        `ifdef SRAM_IP
        .INSTANTIATE_ASIC_MEMORY(1'b1),
        `else
        .INSTANTIATE_ASIC_MEMORY(1'b0),
        `endif
        .INIT_MEMORY_ON_RESET('0) // HPDC doesn't initialize any SRAM
    ) sram (
        `ifdef INTEL_PHYSICAL_MEM_CTRL
        .INTEL_MEM_CTRL(uhdusplr_mem_ctrl),
        `endif
        .SR_ID('0),
        .clk(clk),
        .rst_n(rst_n),
        .clk_en(cs),
        .rdw_en(we),
        .addr(addr),
        .data_in(wdata),
        .data_mask_in({DATA_SIZE{we}}),
        .data_out(rdata),
        .srams_rtap_data( /* Unconnected */ ),
        .rtap_srams_bist_command('0),
        .rtap_srams_bist_data('0)
    );

endmodule : hpdcache_sram
